LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
ENTITY Calculator IS

PORT 
(
CLOCK_50 : IN STD_LOGIC;	
KEY : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
DRAM_CLK, DRAM_CKE : OUT STD_LOGIC;
DRAM_ADDR : OUT STD_LOGIC_VECTOR(11 DOWNTO 0);
DRAM_BA_1, DRAM_BA_0 : BUFFER STD_LOGIC;
DRAM_CS_N, DRAM_CAS_N, DRAM_RAS_N, DRAM_WE_N : OUT STD_LOGIC;
DRAM_DQ : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
DRAM_UDQM, DRAM_LDQM : BUFFER STD_LOGIC;
LEDG   : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
LCD_EN : OUT STD_LOGIC;
LCD_RW : OUT STD_LOGIC;
LCD_RS : OUT STD_LOGIC;
LCD_ON : OUT STD_LOGIC;
LCD_DATA : INOUT STD_LOGIC_VECTOR(7 DOWNTO 0)
);
END Calculator;

ARCHITECTURE Structure OF Calculator IS
COMPONENT nios_system
PORT ( 
              -- 1) global signals:
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- the_LCD
                 signal LCD_E_from_the_LCD : OUT STD_LOGIC;
                 signal LCD_RS_from_the_LCD : OUT STD_LOGIC;
                 signal LCD_RW_from_the_LCD : OUT STD_LOGIC;
                 signal LCD_data_to_and_from_the_LCD : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0);

              -- the_sdram
                 signal zs_addr_from_the_sdram : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
                 signal zs_ba_from_the_sdram : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal zs_cas_n_from_the_sdram : OUT STD_LOGIC;
                 signal zs_cke_from_the_sdram : OUT STD_LOGIC;
                 signal zs_cs_n_from_the_sdram : OUT STD_LOGIC;
                 signal zs_dq_to_and_from_the_sdram : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal zs_dqm_from_the_sdram : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal zs_ras_n_from_the_sdram : OUT STD_LOGIC;
                 signal zs_we_n_from_the_sdram : OUT STD_LOGIC
      );

END COMPONENT;

COMPONENT sdram_pll
PORT ( 
		inclk0 	: IN STD_LOGIC;
		c0 		: OUT STD_LOGIC );
END COMPONENT;

SIGNAL BA : STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL DQM : STD_LOGIC_VECTOR(1 DOWNTO 0);

BEGIN

-- Instantiate the Nios II system entity generated by the SOPC Builder.
NiosII: nios_system 
PORT MAP 
(
--Global mappings
clk => CLOCK_50, 
reset_n => KEY(0), 
--LCD mappings
LCD_E_from_the_LCD => LCD_EN,
LCD_RS_from_the_LCD => LCD_RS,
LCD_RW_from_the_LCD => LCD_RW,
LCD_data_to_and_from_the_LCD => LCD_DATA, 
--SDRAM mappings
zs_addr_from_the_sdram => DRAM_ADDR, 
zs_ba_from_the_sdram => BA, 
zs_cas_n_from_the_sdram => DRAM_CAS_N, 
zs_cke_from_the_sdram => DRAM_CKE, 
zs_cs_n_from_the_sdram => DRAM_CS_N,
zs_dq_to_and_from_the_sdram => DRAM_DQ, 
zs_dqm_from_the_sdram => DQM, 
zs_ras_n_from_the_sdram => DRAM_RAS_N, 
zs_we_n_from_the_sdram =>DRAM_WE_N 
);

-- Instantiate the entity sdram_pll (inclk0, c0).
neg_3ns: sdram_pll 
PORT MAP
(
inclk0 => CLOCK_50, 
c0 => DRAM_CLK
);

LCD_ON <= '1';

DRAM_BA_1 <= BA(1);
DRAM_BA_0 <= BA(0);

DRAM_UDQM <= DQM(1);
DRAM_LDQM <= DQM(0);
	
END Structure;